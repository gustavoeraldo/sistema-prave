* C:\Users\Gustavo\Downloads\UFRN2SEASON\emg_pspice\instrumetation_amp.sch

* Schematics Version 9.1 - Web Update 1
* Fri Mar 12 12:17:50 2021



** Analysis setup **
.tran 0ns 50ms 0 1m
.OP 
.STMLIB "emg2.stl"


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "instrumetation_amp.net"
.INC "instrumetation_amp.als"


.probe


.END
