* C:\Users\Gustavo\Downloads\UFRN2SEASON\emg_pspice\emg_circut.sch

* Schematics Version 9.1 - Web Update 1
* Fri Mar 12 23:46:37 2021



** Analysis setup **
.tran 0ns 80ms 0 1ms
.OP 
.STMLIB "emg_circut.stl"


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "emg_circut.net"
.INC "emg_circut.als"


.probe


.END
